module state_update#(
	parameter N = 32,
	parameter Q = 18,
	parameter T = 0.00001
)
(	input signed [N-1:0] ialpha,ibeta,omega,theta,
	input clk,reset,
	output signed [N-1:0] ialphae,ibetae,omegae,thetae
	);



endmodule